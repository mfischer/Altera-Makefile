module top_level (input CLOCK_50);

// This is a template

endmodule
